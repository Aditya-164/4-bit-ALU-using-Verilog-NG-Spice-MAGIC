* SPICE3 file created from AND3.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)

M1000 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=95 ps=78
M1001 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=86 ps=52
M1002 not_0/in C a_2_n39# Gnd CMOSN w=6 l=2
+  ad=84 pd=40 as=114 ps=50
M1003 not_0/in C vdd w_n31_n3# CMOSP w=5 l=2
+  ad=90 pd=66 as=0 ps=0
M1004 not_0/in A vdd w_n31_n3# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_2_n39# B a_n18_n39# Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=108 ps=48
M1006 not_0/in B vdd w_n31_n3# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_n18_n39# A gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n31_n3# C 0.08fF
C1 vdd w_n31_n3# 0.14fF
C2 out gnd 0.08fF
C3 not_0/in out 0.02fF
C4 not_0/w_n9_1# not_0/in 0.06fF
C5 w_n31_n3# B 0.08fF
C6 not_0/in C 0.12fF
C7 not_0/in w_n31_n3# 0.10fF
C8 not_0/in vdd 0.24fF
C9 not_0/w_n9_1# out 0.03fF
C10 w_n31_n3# A 0.08fF
C11 not_0/in B 0.12fF
C12 not_0/in gnd 0.01fF
C13 vdd out 0.07fF
C14 not_0/w_n9_1# vdd 0.05fF
C15 C Gnd 0.29fF
C16 B Gnd 0.28fF
C17 A Gnd 0.29fF
C18 w_n31_n3# Gnd 0.80fF
C19 gnd Gnd 0.24fF
C20 out Gnd 0.11fF
C21 vdd Gnd 0.16fF
C22 not_0/in Gnd 0.26fF
C23 not_0/w_n9_1# Gnd 0.40fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(C)+4 v(Out)+6

.end
.endc

