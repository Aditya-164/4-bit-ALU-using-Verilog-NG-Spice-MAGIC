* SPICE3 file created from OR4.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)
V_in_d D gnd PULSE(0 1.8 0ns 100ps 100ps 120ns 150ns)

M1000 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=45 ps=38
M1001 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=188 ps=122
M1002 not_0/in A gnd Gnd CMOSN w=6 l=2
+  ad=150 pd=98 as=0 ps=0
M1003 not_0/in D gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_30_9# C a_10_9# w_n21_0# CMOSP w=5 l=2
+  ad=90 pd=46 as=90 ps=46
M1005 a_n8_9# A vdd w_n21_0# CMOSP w=5 l=2
+  ad=80 pd=42 as=0 ps=0
M1006 a_10_9# B a_n8_9# w_n21_0# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 not_0/in D a_30_9# w_n21_0# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1008 not_0/in B gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 not_0/in C gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 not_0/w_n9_1# vdd 0.05fF
C1 not_0/in D 0.09fF
C2 w_n21_0# B 0.08fF
C3 C not_0/in 0.06fF
C4 out not_0/in 0.02fF
C5 w_n21_0# not_0/in 0.04fF
C6 not_0/w_n9_1# not_0/in 0.06fF
C7 not_0/in vdd 0.02fF
C8 out gnd 0.08fF
C9 w_n21_0# A 0.08fF
C10 B not_0/in 0.06fF
C11 w_n21_0# D 0.09fF
C12 w_n21_0# C 0.08fF
C13 out not_0/w_n9_1# 0.03fF
C14 gnd not_0/in 0.45fF
C15 out vdd 0.07fF
C16 w_n21_0# vdd 0.11fF
C17 D Gnd 0.34fF
C18 C Gnd 0.35fF
C19 B Gnd 0.20fF
C20 A Gnd 0.20fF
C21 w_n21_0# Gnd 1.84fF
C22 gnd Gnd 0.74fF
C23 out Gnd 0.11fF
C24 vdd Gnd 0.25fF
C25 not_0/in Gnd 0.69fF
C26 not_0/w_n9_1# Gnd 0.40fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(C)+4 v(D)+6 v(Out)+8

.end
.endc
