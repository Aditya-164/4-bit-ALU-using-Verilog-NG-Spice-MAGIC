* SPICE3 file created from AND4.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)
V_in_d D gnd PULSE(0 1.8 0ns 100ps 100ps 90ns 130ns)


M1000 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=135 ps=104
M1001 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=60 ps=44
M1002 a_25_n36# C a_6_n36# Gnd CMOSN w=5 l=2
+  ad=85 pd=44 as=85 ps=44
M1003 not_0/in B vdd w_n27_2# CMOSP w=5 l=2
+  ad=105 pd=82 as=0 ps=0
M1004 not_0/in C vdd w_n27_2# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 not_0/in A vdd w_n27_2# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 not_0/in D vdd w_n27_2# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 not_0/in D a_25_n36# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 a_6_n36# B a_n14_n36# Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=90 ps=46
M1009 a_n14_n36# A gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 not_0/in not_0/w_n9_1# 0.06fF
C1 not_0/in gnd 0.05fF
C2 not_0/in out 0.02fF
C3 C not_0/in 0.06fF
C4 vdd not_0/w_n9_1# 0.05fF
C5 w_n27_2# not_0/in 0.13fF
C6 w_n27_2# B 0.08fF
C7 vdd out 0.07fF
C8 w_n27_2# vdd 0.18fF
C9 not_0/in B 0.06fF
C10 out not_0/w_n9_1# 0.03fF
C11 w_n27_2# D 0.08fF
C12 gnd out 0.08fF
C13 vdd not_0/in 0.38fF
C14 w_n27_2# C 0.08fF
C15 not_0/in D 0.06fF
C16 A w_n27_2# 0.08fF
C17 D Gnd 0.31fF
C18 C Gnd 0.31fF
C19 B Gnd 0.30fF
C20 A Gnd 0.29fF
C21 w_n27_2# Gnd 1.58fF
C22 gnd Gnd 0.28fF
C23 out Gnd 0.10fF
C24 vdd Gnd 0.30fF
C25 not_0/in Gnd 0.31fF
C26 not_0/w_n9_1# Gnd 0.40fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(C)+4 v(D)+6 v(Out)+8

.end
.endc

