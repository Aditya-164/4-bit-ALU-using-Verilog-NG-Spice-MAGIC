* SPICE3 file created from OR3.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)


M1000 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=62 ps=44
M1001 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=224 ps=122
M1002 not_0/in C gnd Gnd CMOSN w=6 l=2
+  ad=186 pd=98 as=0 ps=0
M1003 a_n42_10# A vdd w_n59_4# CMOSP w=6 l=2
+  ad=150 pd=62 as=0 ps=0
M1004 a_n15_10# B a_n42_10# w_n59_4# CMOSP w=6 l=2
+  ad=186 pd=74 as=0 ps=0
M1005 not_0/in A gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 not_0/in B gnd Gnd CMOSN w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 not_0/in C a_n15_10# w_n59_4# CMOSP w=6 l=2
+  ad=90 pd=42 as=0 ps=0
C0 w_n59_4# C 0.06fF
C1 vdd w_n59_4# 0.15fF
C2 out gnd 0.08fF
C3 not_0/in out 0.02fF
C4 not_0/w_n9_1# not_0/in 0.06fF
C5 w_n59_4# B 0.06fF
C6 not_0/in C 0.08fF
C7 not_0/in w_n59_4# 0.03fF
C8 not_0/in vdd 0.02fF
C9 not_0/w_n9_1# out 0.03fF
C10 w_n59_4# A 0.06fF
C11 not_0/in B 0.08fF
C12 not_0/in gnd 0.06fF
C13 vdd out 0.07fF
C14 not_0/w_n9_1# vdd 0.05fF
C15 C Gnd 0.74fF
C16 B Gnd 0.11fF
C17 A Gnd 0.76fF
C18 w_n59_4# Gnd 2.25fF
C19 gnd Gnd 0.99fF
C20 out Gnd 0.11fF
C21 vdd Gnd 0.88fF
C22 not_0/in Gnd 1.13fF
C23 not_0/w_n9_1# Gnd 0.40fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(C)+4 v(Out)+6

.end
.endc
