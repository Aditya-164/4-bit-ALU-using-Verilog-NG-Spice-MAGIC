* SPICE3 file created from AND.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

M1000 not_0/in B vdd NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=40 pd=36 as=68 ps=58
M1001 not_0/in B NAND_0/a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1002 not_0/in A vdd NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 NAND_0/a_13_n30# A gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=80 ps=52
M1004 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 out not_0/w_n9_1# 0.03fF
C1 out not_0/in 0.02fF
C2 A B 0.02fF
C3 vdd not_0/w_n9_1# 0.05fF
C4 gnd not_0/in 0.01fF
C5 vdd not_0/in 0.21fF
C6 B not_0/in 0.09fF
C7 not_0/w_n9_1# not_0/in 0.06fF
C8 A NAND_0/w_n1_n1# 0.06fF
C9 vdd NAND_0/w_n1_n1# 0.09fF
C10 B NAND_0/w_n1_n1# 0.06fF
C11 NAND_0/w_n1_n1# not_0/in 0.07fF
C12 out gnd 0.08fF
C13 out vdd 0.07fF
C14 gnd Gnd 1.19fF
C15 out Gnd 0.08fF
C16 vdd Gnd 1.80fF
C17 not_0/in Gnd 0.43fF
C18 not_0/w_n9_1# Gnd 0.40fF
C19 B Gnd 0.27fF
C20 A Gnd 0.27fF
C21 NAND_0/w_n1_n1# Gnd 0.69fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(Out)+4

.end
.endc
