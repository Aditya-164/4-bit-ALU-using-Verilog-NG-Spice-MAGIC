* SPICE3 file created from decoder.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_s0 s0 gnd dc 0
V_in_s1 s1 gnd dc 0

M1000 AND_0/not_0/in AND_1/B vdd AND_0/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=40 pd=36 as=312 ps=268
M1001 AND_0/not_0/in AND_1/B AND_0/NAND_0/a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1002 AND_0/not_0/in AND_2/B vdd AND_0/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 AND_0/NAND_0/a_13_n30# AND_2/B gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=360 ps=244
M1004 en0 AND_0/not_0/in vdd AND_0/not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 en0 AND_0/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1006 AND_1/not_0/in AND_1/B vdd AND_1/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1007 AND_1/not_0/in AND_1/B AND_1/NAND_0/a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1008 AND_1/not_0/in s0 vdd AND_1/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 AND_1/NAND_0/a_13_n30# s0 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 en1 AND_1/not_0/in vdd AND_1/not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 en1 AND_1/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1012 AND_2/not_0/in AND_2/B vdd AND_2/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1013 AND_2/not_0/in AND_2/B AND_2/NAND_0/a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1014 AND_2/not_0/in s1 vdd AND_2/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 AND_2/NAND_0/a_13_n30# s1 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 en2 AND_2/not_0/in vdd AND_2/not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 en2 AND_2/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 AND_3/not_0/in s0 vdd AND_3/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1019 AND_3/not_0/in s0 AND_3/NAND_0/a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1020 AND_3/not_0/in s1 vdd AND_3/NAND_0/w_n1_n1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 AND_3/NAND_0/a_13_n30# s1 gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 en3 AND_3/not_0/in vdd AND_3/not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1023 en3 AND_3/not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1024 AND_2/B s0 vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1025 AND_2/B s0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1026 AND_1/B s1 vdd not_1/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 AND_1/B s1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 AND_1/B s0 0.52fF
C1 gnd en0 0.08fF
C2 en2 AND_2/not_0/w_n9_1# 0.03fF
C3 AND_0/not_0/w_n9_1# en0 0.03fF
C4 gnd AND_2/B 0.21fF
C5 gnd s0 0.34fF
C6 s0 AND_1/NAND_0/w_n1_n1# 0.06fF
C7 vdd AND_0/NAND_0/w_n1_n1# 0.09fF
C8 vdd AND_3/not_0/w_n9_1# 0.05fF
C9 AND_3/NAND_0/w_n1_n1# s0 0.06fF
C10 not_1/w_n9_1# vdd 0.05fF
C11 en2 gnd 0.08fF
C12 vdd not_0/w_n9_1# 0.05fF
C13 AND_3/not_0/in AND_3/not_0/w_n9_1# 0.06fF
C14 AND_2/not_0/in vdd 0.21fF
C15 gnd AND_1/B 0.33fF
C16 AND_1/B AND_1/NAND_0/w_n1_n1# 0.06fF
C17 AND_0/not_0/in en0 0.02fF
C18 AND_2/B AND_2/NAND_0/w_n1_n1# 0.06fF
C19 vdd en1 0.15fF
C20 vdd AND_3/not_0/in 0.21fF
C21 s1 AND_2/B 1.25fF
C22 s1 s0 0.85fF
C23 AND_0/NAND_0/w_n1_n1# AND_2/B 0.06fF
C24 en3 gnd 0.08fF
C25 vdd AND_1/not_0/w_n9_1# 0.05fF
C26 vdd AND_1/not_0/in 0.21fF
C27 AND_1/B AND_0/not_0/in 0.09fF
C28 en1 AND_1/not_0/w_n9_1# 0.03fF
C29 AND_2/B not_0/w_n9_1# 0.03fF
C30 s1 AND_1/B 0.02fF
C31 en1 AND_1/not_0/in 0.02fF
C32 AND_2/not_0/in AND_2/B 0.09fF
C33 s0 not_0/w_n9_1# 0.06fF
C34 vdd en0 0.15fF
C35 gnd AND_0/not_0/in 0.01fF
C36 vdd AND_2/B 0.15fF
C37 AND_0/not_0/in AND_0/not_0/w_n9_1# 0.06fF
C38 AND_0/NAND_0/w_n1_n1# AND_1/B 0.06fF
C39 vdd s0 0.10fF
C40 s1 gnd 0.45fF
C41 AND_2/not_0/in en2 0.02fF
C42 not_1/w_n9_1# AND_1/B 0.03fF
C43 s1 AND_3/NAND_0/w_n1_n1# 0.06fF
C44 en2 vdd 0.15fF
C45 AND_1/not_0/w_n9_1# AND_1/not_0/in 0.06fF
C46 AND_2/not_0/in AND_2/not_0/w_n9_1# 0.06fF
C47 AND_3/not_0/in s0 0.09fF
C48 AND_2/not_0/w_n9_1# vdd 0.05fF
C49 vdd AND_1/B 0.07fF
C50 AND_2/not_0/in gnd 0.01fF
C51 en3 AND_3/not_0/w_n9_1# 0.03fF
C52 vdd AND_1/NAND_0/w_n1_n1# 0.09fF
C53 vdd AND_0/not_0/w_n9_1# 0.05fF
C54 s1 AND_2/NAND_0/w_n1_n1# 0.06fF
C55 AND_3/NAND_0/w_n1_n1# vdd 0.09fF
C56 en1 gnd 0.08fF
C57 AND_2/B s0 0.21fF
C58 AND_0/NAND_0/w_n1_n1# AND_0/not_0/in 0.07fF
C59 AND_3/not_0/in gnd 0.01fF
C60 vdd en3 0.07fF
C61 AND_1/B AND_1/not_0/in 0.09fF
C62 AND_3/NAND_0/w_n1_n1# AND_3/not_0/in 0.07fF
C63 not_1/w_n9_1# s1 0.06fF
C64 AND_2/not_0/in AND_2/NAND_0/w_n1_n1# 0.07fF
C65 gnd AND_1/not_0/in 0.01fF
C66 AND_1/NAND_0/w_n1_n1# AND_1/not_0/in 0.07fF
C67 vdd AND_2/NAND_0/w_n1_n1# 0.09fF
C68 en3 AND_3/not_0/in 0.02fF
C69 AND_2/B AND_1/B 0.41fF
C70 vdd AND_0/not_0/in 0.21fF
C71 not_1/w_n9_1# Gnd 0.40fF
C72 not_0/w_n9_1# Gnd 0.40fF
C73 en3 Gnd 0.15fF
C74 AND_3/not_0/w_n9_1# Gnd 0.40fF
C75 gnd Gnd 22.68fF
C76 AND_3/not_0/in Gnd 0.43fF
C77 vdd Gnd 7.36fF
C78 s0 Gnd 7.82fF
C79 s1 Gnd 3.71fF
C80 AND_3/NAND_0/w_n1_n1# Gnd 0.69fF
C81 en2 Gnd 0.18fF
C82 AND_2/not_0/w_n9_1# Gnd 0.40fF
C83 AND_2/not_0/in Gnd 0.43fF
C84 AND_2/B Gnd 0.69fF
C85 AND_2/NAND_0/w_n1_n1# Gnd 0.69fF
C86 AND_1/not_0/w_n9_1# Gnd 0.40fF
C87 AND_1/not_0/in Gnd 0.43fF
C88 AND_1/B Gnd 0.69fF
C89 AND_1/NAND_0/w_n1_n1# Gnd 0.69fF
C90 en0 Gnd 0.15fF
C91 AND_0/not_0/w_n9_1# Gnd 0.40fF
C92 AND_0/not_0/in Gnd 0.43fF
C93 AND_0/NAND_0/w_n1_n1# Gnd 0.69fF


.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(s0) v(s1)+2 v(en0)+4 v(en1)+6 v(en2)+8 v(en3)+10 

.end
.endc
