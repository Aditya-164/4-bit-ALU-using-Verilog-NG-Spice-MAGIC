* SPICE3 file created from AND5.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 100ns)
V_in_d D gnd PULSE(0 1.8 0ns 100ps 100ps 90ns 130ns)
V_in_e E gnd PULSE(0 1.8 0ns 100ps 100ps 120ns 160ns)

M1000 out not_0/in vdd not_0/w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=155 ps=122
M1001 out not_0/in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=52 ps=42
M1002 a_10_n35# B a_n9_n35# Gnd CMOSN w=4 l=2
+  ad=68 pd=42 as=68 ps=42
M1003 not_0/in E vdd w_n22_7# CMOSP w=5 l=2
+  ad=140 pd=106 as=0 ps=0
M1004 not_0/in B vdd w_n22_7# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 not_0/in C vdd w_n22_7# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_29_n35# C a_10_n35# Gnd CMOSN w=4 l=2
+  ad=72 pd=44 as=0 ps=0
M1007 not_0/in E a_49_n35# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=68 ps=42
M1008 a_n9_n35# A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_49_n35# D a_29_n35# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 not_0/in D vdd w_n22_7# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 not_0/in A vdd w_n22_7# CMOSP w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 not_0/in B 0.06fF
C1 A w_n22_7# 0.08fF
C2 vdd not_0/w_n9_1# 0.05fF
C3 out not_0/w_n9_1# 0.03fF
C4 w_n22_7# not_0/in 0.17fF
C5 w_n22_7# B 0.08fF
C6 gnd out 0.08fF
C7 vdd out 0.07fF
C8 not_0/in D 0.06fF
C9 w_n22_7# D 0.08fF
C10 not_0/in not_0/w_n9_1# 0.06fF
C11 not_0/in gnd 0.03fF
C12 vdd not_0/in 0.34fF
C13 not_0/in out 0.02fF
C14 C not_0/in 0.06fF
C15 w_n22_7# vdd 0.26fF
C16 w_n22_7# C 0.08fF
C17 not_0/in E 0.09fF
C18 w_n22_7# E 0.08fF
C19 E Gnd 0.32fF
C20 D Gnd 0.32fF
C21 C Gnd 0.32fF
C22 B Gnd 0.32fF
C23 A Gnd 0.32fF
C24 w_n22_7# Gnd 2.15fF
C25 gnd Gnd 0.32fF
C26 out Gnd 0.11fF
C27 vdd Gnd 0.47fF
C28 not_0/in Gnd 0.36fF
C29 not_0/w_n9_1# Gnd 0.40fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(C)+4 v(D)+6 v(E)+8 v(Out)+10

.end
.endc

