.include TSMC_180nm.txt
.include fulladder.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c C gnd dc 'SUPPLY'

X1 A B C S Car vdd gnd fulladder

* X1 node_a node_b node_c node_x gnd NAND
* X2 node_a node_c node_d node_x gnd NAND
* X3 node_b node_c node_e node_x gnd NAND
* X4 node_e node_d node_out node_x gnd NAND


C1 S gnd 100f
C2 Car gnd 100f

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(A) v(B)+2 v(C)+4 v(S)+6 v(Car)+8
hardcopy image.ps v(A) v(B)+2 v(C)+4 v(S)+6 v(Car)+8
.end
.endc