* SPICE3 file created from NAND.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

M1000 out B vdd vdd# CMOSP w=4 l=2
+  ad=40 pd=36 as=48 ps=40
M1001 out B a_13_n30# Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=80 ps=42
M1002 out A vdd vdd# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_13_n30# A gnd Gnd CMOSN w=5 l=2
+  ad=0 pd=0 as=60 ps=34
C0 out vdd 0.21fF
C1 vdd# A 0.06fF
C2 vdd# B 0.06fF
C3 vdd# vdd 0.09fF
C4 vdd# out 0.07fF
C5 out B 0.09fF

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(A) v(B)+2 v(Out)+4

.end
.endc
